// SRAM 高速缓存
module  SRAM(input a,b,output  out);
	



endmodule;
