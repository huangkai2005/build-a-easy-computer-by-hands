module SRFF (input R, clock, S, output Q, Q_dot);
  // your code here

endmodule

