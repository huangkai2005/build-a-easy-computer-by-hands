
module HalfAdder(input a,b, output sum, carry);
  // your code here

endmodule

