
module Not(input in, output out);
  // your code here
	nand n(out,in,in);
endmodule



