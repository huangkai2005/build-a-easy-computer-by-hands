

module RAM512(input [15:0] in, input clk,load, input [8:0] address, output [15:0] out);
    // your code here

endmodule
