module DFF(input in, clock, load, output out);
  // your code here

endmodule

