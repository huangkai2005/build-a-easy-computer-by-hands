module IsNeg(input[15:0] in, output out);
  // your code here

endmodule
