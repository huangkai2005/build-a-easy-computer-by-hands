
module Not(input in, output out);
  // your code here

endmodule



