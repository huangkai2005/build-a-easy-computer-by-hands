module IsNeg(input[15:0] in, output out);
  // your code here
	and a(out,in[15],1);
endmodule
