
module Or(input a, b, output out);
  // your code here

endmodule
