/**
 * 16-way Or: 
 * out = (in[0] or in[1] or ... or in[15])
 */

module Or16Way(input[15:0] in,output out);
    // your code here

endmodule


